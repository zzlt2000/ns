module loss (
    input   signed  wire    [NTOTAL_BITS-1:0] rays_count;
    input   [8:0]valid;     //输出信号
);
    
endmodule